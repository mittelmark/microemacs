// -!- v-lang -!-
module main

pub fn test () {
    
}

fn main() {
    println("Hello V World!")
}
